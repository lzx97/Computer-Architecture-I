// Test bench for ALU
`timescale 1ns/10ps

// Meaning of signals in and out of the ALU:

// Flags:
// negative: whether the result output is negative if interpreted as 2's comp.
// zero: whether the result output was a 64-bit zero.
// overflow: on an add or subtract, whether the computation overflowed if the inputs are interpreted as 2's comp.
// carry_out: on an add or subtract, whether the computation produced a carry-out.

// cntrl			Operation						Notes:
// 000:			result = B					value of overflow and carry_out unimportant
// 001			result = A (<< or >>) B		value of overflow and carry_out unimportant
// 010:			result = A + B
// 011:			result = A - B
// 100:			result = bitwise A & B		value of overflow and carry_out unimportant
// 101:			result = bitwise A | B		value of overflow and carry_out unimportant
// 110:			result = bitwise A XOR B	value of overflow and carry_out unimportant
// 111:			result = A * B				value of overflow and carry_out unimportant

module alustim();

	parameter delay = 100000;

	logic		[63:0]	A, B;
	logic		[2:0]		cntrl;
	logic 				shiftdir;
	logic		[63:0]	result;
	logic					negative, zero, overflow, carry_out;

	parameter ALU_PASS_B=3'b000, ALU_ADD=3'b010, ALU_SUBTRACT=3'b011, ALU_AND=3'b100, ALU_OR=3'b101, ALU_XOR=3'b110, ALU_SHIFT=3'b001, ALU_MUL= 3'b111;
	

	alu dut (.A, .B, .cntrl, .result, .negative, .zero, .overflow, .carry_out, .shiftdir);

	// Force %t's to print in a nice format.
	initial $timeformat(-9, 2, " ns", 10);

	integer i;
	logic [63:0] test_val;
	initial begin
	
		$display("%t testing PASS_B operations", $time);
		cntrl = ALU_PASS_B;
		for (i=0; i<100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == B && negative == B[63] && zero == (B == 0));
		end
		
		$display("%t testing addition", $time);
		cntrl = ALU_ADD;
			for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A + B) && negative == result[63] && zero == (result == 0) && overflow == ((~A[63] & ~B[63] & result[63]) | (A[63] & B[63] & ~result[63])));
		end
		A = 64'h0000000000000001; B = 64'h0000000000000001;
		#(delay);
		assert(result == 64'h0000000000000002 && carry_out == 0 && overflow == 0 && negative == 0 && zero == 0);
		
		A = 64'h7fffffffffffffff; B = 64'h1;
		#(delay);
		assert(result == 64'h8000000000000000 && carry_out == 0 && overflow == 1 && negative == 1 && zero == 0);
		
		A = 64'h8000000000000000; B = 64'h8000000000000000;
		#(delay);
		assert(result == 64'h0000000000000000 && carry_out == 1 && overflow == 1 && negative == 0 && zero == 1);
		
		
		$display("%t testing subtraction", $time);
		cntrl = ALU_SUBTRACT;
		for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A - B) && negative == result[63] && zero == (result == 0) && overflow == ((~A[63] & B[63] & result[63]) | (A[63] & ~B[63] & ~result[63])));
		end

		A = 64'h1; B = 64'h2;
		#(delay);
		assert(result == 64'hffffffffffffffff && carry_out == 0 && overflow == 0 && negative == 1 && zero == 0);
		
		A = 64'h7fffffffffffffff; B = 64'hffffffffffffffff;
		#(delay);
		assert(result == 64'h8000000000000000 && carry_out == 0 && overflow == 1 && negative == 1 && zero == 0);
		
		A = 100; B = 10000;
		#(delay);
		assert(result == -9900);
		
		$display("%t testing and", $time);
		cntrl = ALU_AND;
		for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A & B) && negative == result[63] && zero == (result == 0));
		end
		
		
		$display("%t testing or", $time);
		cntrl = ALU_OR;
		for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A | B) && negative == result[63] && zero == (result == 0));
		end
		
		$display("%t testing xor", $time);
		cntrl = ALU_XOR;
		for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A ^ B) && negative == result[63] && zero == (result == 0));
		end

		$display("%t testing shift", $time);
		cntrl = ALU_SHIFT;
		shiftdir = 0;
		for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A << B[5:0]));
		end

		shiftdir = 1;
		for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A >> B[5:0]));
		end

		$display("%t testing multiply", $time);
		cntrl = ALU_MUL;
		for (i = 0; i < 100; i++) begin
			A = $random(); B = $random();
			#(delay);
			assert(result == (A * B));
		end
	end
endmodule 