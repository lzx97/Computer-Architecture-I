module forwaring();
	input [4:0] Rn, Rd;
	input [4:0] Rd_EX_MEM, Rd_MEM_WBl;
	input [] cntrl_EX_MEM, cntrl_MEM_WB; // fix width?
	output [1:0] muxcntrl0, muxcntrl1;
	

endmodule 